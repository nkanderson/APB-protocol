// FIXME: This file is a placeholder for testing project directory setup
// and compilation scripting. Modify, edit, or delete this file as necessary
// once development begins.
package apb_pkg;
// Add basic typedefs, parameters, etc.
endpackage
